module mkPPP(MessageGet c2m, MessagePut m2c, WideMem mem, Empty ifc);

endmodule
